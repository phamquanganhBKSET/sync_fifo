`define FIFO_DEPTH 256
`define DATA_WIDTH 32
`define FIFO_DEPTH 8
`define DATA_WIDTH 32